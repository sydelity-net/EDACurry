Alter command example
r1 1 2 1k
r2 2 0 1k
c1 2 0 1n
.ac dec 10 200 1000meg
vin 1 0 ac 1

.plot ac vdb(2) (-90, 0)

.alter
    r1 1 2 10k
    c1 2 0 100p
    .ac dec 15 200 1500meg
.end

.param RVAL=1k
.param MULT=1
.alter first
    .param RVAL=1.3k
    .param MULT=1.3
.alter second
    .param RVAL=0.7k
    .param MULT=1.3
.alter
    .param RVAL=0.7k
    .param MULT=0.7
.alter fourth
    .param RVAL=1.3k
    .param MULT=0.7
.end

r1 1 0 1
r2 2 0 1
.alter 1
r1 1 0 2
.alter 2
r2 2 0 2
