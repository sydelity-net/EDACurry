// ============================================================================
// SPICE
// ============================================================================
.tran 2e-6 2e-3