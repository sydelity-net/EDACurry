// ============================================================================
// SPICE
// ============================================================================
*Model for NMOS Transistor
.MODEL nfet NMOS ( LEVEL = 8
    +VERSION = 3.2 TNOM = 27 TOX = 1.42E-8
    +NCH = 1.7E17 VTH0 = 0.6106006
    +K1 = 0.8791418 K2 = -0.0928691 K3 = 18.3613087
    +K3B = -8.1787847 W0 = 1E-8 NLX = 1E-9
    +DVT0W = 0 DVT1W = 0 DVT2W = 0
    +DVT0 = 3.5655768 DVT1 = 0.3802648 DVT2 = -0.0874051
    +U0 = 452.6968866 UA = 1.406301E-13 UB = 1.618501E-18
    +UC = 5.36169E-12 VSAT = 1.802287E5 A0 = 0.5750334
    +AGS = 0.1061895 B0 = 2.728576E-6 B1 = 5E-6
    +KETA = -8.123787E-5 A1 = 4.190554E-4 A2 = 0.3323258
    +RDSW = 1.06188E3 PRWG = 0.0883334 PRWB = 0.0315574
    +WR = 1 WINT = 2.308608E-7 LINT = 7.347987E-8
    +XL = 1E-7 DWG = -1.605516E-8
    +DWB = 3.927415E-8 VOFF = 0 NFACTOR = 0.4571776
    +CIT = 0 CDSC = 2.4E-4 CDSCD = 0
    +CDSCB = 0 ETA0 = 2.176689E-3 ETAB = -8.669487E-5
    +DSUB = 0.0553447 PCLM = 2.4898877 PDIBLC1 = 1
    +PDIBLC2 = 2.156583E-3 PDIBLCB = -0.0394428 DROUT = 0.9016259
    +PSCBE1 = 6.238215E8 PSCBE2 = 1.760403E-4 PVAG = 0
    +DELTA = 0.01 RSH = 83.8 MOBMOD = 1
    +PRT = 0 UTE = -1.5 KT1 = -0.11
    +KT1L = 0 KT2 = 0.022 UA1 = 4.31E-9
    +UB1 = -7.61E-18 UC1 = -5.6E-11 AT = 3.3E4
    +WL = 0 WLN = 1 WW = 0
    +WWN = 1 WWL = 0 LL = 0
    +LLN = 1 LW = 0 LWN = 1
    +LWL = 0 CAPMOD = 2 XPART = 0.5
    +CGDO = 1.97E-10 CGSO = 1.97E-10 CGBO = 1E-9
    +CJ = 4.315315E-4 PB = 0.9194059 MJ = 0.4344423
    +CJSW = 3.335714E-10 PBSW = 0.8 MJSW = 0.1985616
    +CJSWG = 1.64E-10 PBSWG = 0.8 MJSWG = 0.1985616
    +CF = 0 PVTH0 = 0.1570368 PRDSW = 187.3761409
    +PK2 = -0.0254353 WKETA = -0.0181601 LKETA = 1.265053E-3 )

* Model for PMOS Transistor
.MODEL pfet PMOS ( LEVEL = 8
    +VERSION = 3.2 TNOM = 27 TOX = 1.42E-8
    +NCH = 1.7E17 VTH0 = -0.9836276
    +K1 = 0.5265664 K2 = 0.0213923 K3 = 4.4911263
    +K3B = -0.6532905 W0 = 1E-8 NLX = 1E-9
    +DVT0W = 0 DVT1W = 0 DVT2W = 0
    +DVT0 = 2.6487289 DVT1 = 0.4862165 DVT2 = -0.0896609
    +U0 = 222.1424772 UA = 3.307877E-9 UB = 2.667897E-21
    +UC = -5.80948E-11 VSAT = 2E5 A0 = 0.8813584
    +AGS = 0.1156322 B0 = 7.044894E-7 B1 = 3.350124E-6
    +KETA = 4.719307E-4 A1 = 0 A2 = 0.3
    +RDSW = 3E3 PRWG = -0.0562354 PRWB = -5.560433E-3
    +WR = 1 WINT = 2.962387E-7 LINT = 9.667582E-8
    +XL = 1E-7 DWG = -3.741786E-8
    +DWB = 1.377762E-8 VOFF = -0.0788978 NFACTOR = 0.6687895
    +CIT = 0 CDSC = 2.4E-4 CDSCD = 0
    +CDSCB = 0 ETA0 = 0.4372057 ETAB = -0.0880016
    +DSUB = 1 PCLM = 2.1801812 PDIBLC1 = 0.0430345
    +PDIBLC2 = 3.544969E-3 PDIBLCB = -0.0720123 DROUT = 0.2036798
    +PSCBE1 = 5.329158E9 PSCBE2 = 5E-10 PVAG = 0.2660196
    +DELTA = 0.01 RSH = 106.9 MOBMOD = 1
    +PRT = 0 UTE = -1.5 KT1 = -0.11
    +KT1L = 0 KT2 = 0.022 UA1 = 4.31E-9
    +UB1 = -7.61E-18 UC1 = -5.6E-11 AT = 3.3E4
    +WL = 0 WLN = 1 WW = 0
    +WWN = 1 WWL = 0 LL = 0
    +LLN = 1 LW = 0 LWN = 1
    +LWL = 0 CAPMOD = 2 XPART = 0.5
    +CGDO = 2.72E-10 CGSO = 2.72E-10 CGBO = 1E-9
    +CJ = 7.257637E-4 PB = 0.9604987 MJ = 0.4949935
    +CJSW = 3.242689E-10 PBSW = 0.99 MJSW = 0.3345497
    +CJSWG = 6.4E-11 PBSWG = 0.99 MJSWG = 0.3345497
    +CF = 0 PVTH0 = 5.98016E-3 PRDSW = 14.8598424
    +PK2 = 3.73981E-3 WKETA = 3.808346E-3 LKETA = -6.010447E-3 )