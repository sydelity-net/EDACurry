// ============================================================================
// SPICE
// ============================================================================
.tran 2e-6 2e-3

// AC AND TRANSIENT ANALYSIS
.AC    DEC  5    10    10MEG
.TRAN   0.001MS    0.2MS
